Standard cell Simulation
* this file edited to remove everything not in tt lib, makes it a lot faster
.lib "./sky130_fd_pr/models/sky130.lib.spice" tt
* including this file means I can use the cell names without copying them in this file
.include "./sky130_fd_sc_hd.spice"

* 1 inverter
X1_1 A_1  VGND VGND VPWR VPWR Y1_1 sky130_fd_sc_hd__inv_1
C1 Y1_1  VGND 0.1pF

* 2 inverters
X2_1 A_2  VGND VGND VPWR VPWR Y2_1 sky130_fd_sc_hd__inv_1
X2_8 Y2_1 VGND VGND VPWR VPWR Y2_8 sky130_fd_sc_hd__inv_8
C2 Y2_8  VGND 0.1pF

* 3 inverters
X3_1  A_3  VGND VGND VPWR VPWR Y3_1 sky130_fd_sc_hd__inv_1
X3_4  Y3_1 VGND VGND VPWR VPWR Y3_4 sky130_fd_sc_hd__inv_4
X3_16 Y3_4 VGND VGND VPWR VPWR Y3_16 sky130_fd_sc_hd__inv_16
C3 Y3_16 VGND 0.1pF

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create the drive pulse for all 3 chains
Va A_1 VGND pulse(0 1.8 1n 10p 10p 1n 2n)
Vb A_2 VGND pulse(0 1.8 1n 10p 10p 1n 2n)
Vc A_3 VGND pulse(0 1.8 1n 10p 10p 1n 2n)

* setup the transient analysis
.tran 10p 3n 0

.control
run
set color0 = white
set color1 = black
plot A_1 Y1_1 Y2_8 Y3_16
.endc

.end
