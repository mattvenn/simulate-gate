
* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
Va A VGND pulse(0 1.8 1n 10p 10p 1n 2n)
Vb B VGND pulse(0 1.8 1.5n 10p 10p 1n 2n)
.tran 10p 3n 0

.control
run
set color0 = white
set color1 = black
plot A B Y
.endc

.end
